library.ieee;
use iee.std_logic_1164.all;
use iee.numeric_std.all;

entity input_layer is
  port
    (
      
    )
